`include "constants.svh"

module accelerator_tb;
    initial begin
        $display("hello world");
        $finish;
    end
endmodule