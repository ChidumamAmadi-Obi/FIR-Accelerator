`include "constants.v"

`timescale 1ns/1ps

module mac_tb;

endmodule