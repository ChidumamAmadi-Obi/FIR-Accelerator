`include "constants.svh"

module top_tb;
    initial begin
        $display("hello world");  $finish;
    end
endmodule