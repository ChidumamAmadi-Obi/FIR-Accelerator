`include "constants.v"

`timescale 1ns/1ps

module shiftreg_tb;

endmodule