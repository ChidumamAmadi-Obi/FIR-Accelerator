/* TOP WRAPPER TO CONNECT TO THE CV32E40X
*/

`include "constants.svh"
`include "top.sv"

module firAccelerators()

endmodule

