`ifndef CONSTANTS // file guard
`define CONSTANTS

`define DATA_WIDTH 32 // 32 bit mcu
`define NUM_REGS 8

`endif
