`ifndef CONSTANTS // file guard
`define CONSTANTS

`timescale 1ns/1ps
`define DATA_WIDTH 32 // 32 bit mcu
`define NUM_REGS 8

`endif